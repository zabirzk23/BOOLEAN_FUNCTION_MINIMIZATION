library verilog;
use verilog.vl_types.all;
entity Boolean_min_vlg_check_tst is
    port(
        f1              : in     vl_logic;
        f2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Boolean_min_vlg_check_tst;
