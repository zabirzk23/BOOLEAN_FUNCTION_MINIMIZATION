library verilog;
use verilog.vl_types.all;
entity Boolean_min_vlg_vec_tst is
end Boolean_min_vlg_vec_tst;
